`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:09:44 09/04/2017
// Design Name:   testBench
// Module Name:   E:/TE/Winter/VLSI/finalProj/testBench/testBench_tb.v
// Project Name:  testBench
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: testBench
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testBench_tb;
	reg clk;
	reg reset;
	// Outputs
	

	// Instantiate the Unit Under Test (UUT)
	testBench uut (
		
	);

 
	initial begin
		
	end
      
endmodule

